module linter

pub enum IndentStyle {
	tab
	space
	any
}
