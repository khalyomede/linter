module linter

pub struct Linter {
	files []string
	folders []string
	rules Rules
}
