module a

pub fn b() string {
    return "hello world"
}
