module a

fn b() string {
	return "c"
}